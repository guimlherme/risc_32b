library ieee;

use IEEE.STD_LOGIC_1164.ALL;
Use ieee.numeric_std.all ;


entity rom is
	port(
			en			:	in std_logic;
			clk		:	in std_logic;
			Address	:	in std_logic_vector(7 downto 0);
			Data_out:	out std_logic_vector(22 downto 0)
			);
end rom;

architecture rom_a of rom is

type rom is array(0 to 255) of std_logic_vector(22 downto 0);

signal Data_Rom : rom ;



--------------- BEGIN -----------------------------------------------------------------
begin

-- Code here


Data_Rom(0) <= "01100010001000000000000";
Data_Rom(1) <= "01100100000000000000000";
Data_Rom(2) <= "11101000001000110000000";
Data_Rom(3) <= "10100000000000000000000";
Data_Rom(4) <= "11000001011000000000000";
Data_Rom(5) <= "11101000001000100000000";
Data_Rom(6) <= "10100000000000000000000";
Data_Rom(7) <= "11000101001000000000000";
Data_Rom(8) <= "01111010000000000000000";
Data_Rom(9) <= "10100000000000000000000";
Data_Rom(10) <= "11001000000000000000000";
Data_Rom(11) <= "00100010001000000010000";
Data_Rom(12) <= "01001000010000100000000";
Data_Rom(13) <= "10100000000000000000000";
Data_Rom(14) <= "11000011000000000000000";
Data_Rom(15) <= "11101000001000001110000";
Data_Rom(16) <= "10100000000000000000000";
Data_Rom(17) <= "11000011110000000000000";
Data_Rom(18) <= "11101000001000110000000";
Data_Rom(19) <= "10100000000000000000000";
Data_Rom(20) <= "11000001011000000000000";
Data_Rom(21) <= "01111010000000000000000";
Data_Rom(22) <= "10100000000000000000000";
Data_Rom(23) <= "11000000010000000000000";
Data_Rom(24) <= "01001000010000100000000";
Data_Rom(25) <= "10100000000000000000000";
Data_Rom(26) <= "11000011000000000000000";
Data_Rom(27) <= "01111010000000000000000";
Data_Rom(28) <= "10100000000000000000000";
Data_Rom(29) <= "11000001111000000000000";
Data_Rom(30) <= "10001000010000100000000";
Data_Rom(31) <= "10100000000000000000000";
Data_Rom(32) <= "11000100101000000000000";
Data_Rom(33) <= "00000010001000010000000";
Data_Rom(34) <= "01111010000000000000000";
Data_Rom(35) <= "10100000000000000000000";
Data_Rom(36) <= "11000010010000000000000";
Data_Rom(37) <= "00000010001000100000000";
Data_Rom(38) <= "01111010000000000000000";
Data_Rom(39) <= "10100000000000000000000";
Data_Rom(40) <= "11000000010000000000000";
Data_Rom(41) <= "00000010001000000010000";
Data_Rom(42) <= "01001000010000100000000";
Data_Rom(43) <= "10100000000000000000000";
Data_Rom(44) <= "11000110110000000000000";
Data_Rom(45) <= "10001000010000100000000";
Data_Rom(46) <= "10100000000000000000000";
Data_Rom(47) <= "11000111100000000000000";
Data_Rom(48) <= "11101000001000110000000";
Data_Rom(49) <= "10100000000000000000000";
Data_Rom(50) <= "11000000010000000000000";
Data_Rom(51) <= "01111010000000000000000";
Data_Rom(52) <= "10100000000000000000000";
Data_Rom(53) <= "11000101001000000000000";
Data_Rom(54) <= "01001000010000100000000";
Data_Rom(55) <= "10100000000000000000000";
Data_Rom(56) <= "11000110110000000000000";
Data_Rom(57) <= "01111010000000000000000";
Data_Rom(58) <= "10100000000000000000000";
Data_Rom(59) <= "11000101101000000000000";
Data_Rom(60) <= "00100010001000010000000";
Data_Rom(61) <= "01111010000000000000000";
Data_Rom(62) <= "10100000000000000000000";
Data_Rom(63) <= "11000110000000000000000";
Data_Rom(64) <= "10001000010000100000000";
Data_Rom(65) <= "10100000000000000000000";
Data_Rom(66) <= "11001000000000000000000";
Data_Rom(67) <= "00100010001000010000000";
Data_Rom(68) <= "01111010000000000000000";
Data_Rom(69) <= "10100000000000000000000";
Data_Rom(70) <= "11000000010000000000000";





-- Data_Rom(0) <= "01100010001000000000000";
-- Data_Rom(1) <= "01100100000000000000000";
-- Data_Rom(2) <= "11101000001000110000000";
-- Data_Rom(3) <= "11000001110000000000000";
-- Data_Rom(4) <= "10100000000000000000000";
-- Data_Rom(5) <= "10100000000000000000000";
-- Data_Rom(6) <= "11101000001000100000000";
-- Data_Rom(7) <= "11000110101000000000000";
-- Data_Rom(8) <= "10100000000000000000000";
-- Data_Rom(9) <= "10100000000000000000000";
-- Data_Rom(10) <= "01111010000000000000000";
-- Data_Rom(11) <= "11001010011000000000000";
-- Data_Rom(12) <= "10100000000000000000000";
-- Data_Rom(13) <= "10100000000000000000000";
-- Data_Rom(14) <= "00100010001000000010000";
-- Data_Rom(15) <= "01001000010000100000000";
-- Data_Rom(16) <= "11000011111000000000000";
-- Data_Rom(17) <= "10100000000000000000000";
-- Data_Rom(18) <= "10100000000000000000000";
-- Data_Rom(19) <= "11101000001000001110000";
-- Data_Rom(20) <= "11000100111000000000000";
-- Data_Rom(21) <= "10100000000000000000000";
-- Data_Rom(22) <= "10100000000000000000000";
-- Data_Rom(23) <= "11101000001000110000000";
-- Data_Rom(24) <= "11000001110000000000000";
-- Data_Rom(25) <= "10100000000000000000000";
-- Data_Rom(26) <= "10100000000000000000000";
-- Data_Rom(27) <= "01111010000000000000000";
-- Data_Rom(28) <= "11000000010000000000000";
-- Data_Rom(29) <= "10100000000000000000000";
-- Data_Rom(30) <= "10100000000000000000000";
-- Data_Rom(31) <= "01001000010000100000000";
-- Data_Rom(32) <= "11000011111000000000000";
-- Data_Rom(33) <= "10100000000000000000000";
-- Data_Rom(34) <= "10100000000000000000000";
-- Data_Rom(35) <= "01111010000000000000000";
-- Data_Rom(36) <= "11000010011000000000000";
-- Data_Rom(37) <= "10100000000000000000000";
-- Data_Rom(38) <= "10100000000000000000000";
-- Data_Rom(39) <= "10001000010000100000000";
-- Data_Rom(40) <= "11000110000000000000000";
-- Data_Rom(41) <= "10100000000000000000000";
-- Data_Rom(42) <= "10100000000000000000000";
-- Data_Rom(43) <= "00000010001000010000000";
-- Data_Rom(44) <= "01111010000000000000000";
-- Data_Rom(45) <= "11000010111000000000000";
-- Data_Rom(46) <= "10100000000000000000000";
-- Data_Rom(47) <= "10100000000000000000000";
-- Data_Rom(48) <= "00000010001000100000000";
-- Data_Rom(49) <= "01111010000000000000000";
-- Data_Rom(50) <= "11000000010000000000000";
-- Data_Rom(51) <= "10100000000000000000000";
-- Data_Rom(52) <= "10100000000000000000000";
-- Data_Rom(53) <= "00000010001000000010000";
-- Data_Rom(54) <= "01001000010000100000000";
-- Data_Rom(55) <= "11001000110000000000000";
-- Data_Rom(56) <= "10100000000000000000000";
-- Data_Rom(57) <= "10100000000000000000000";
-- Data_Rom(58) <= "10001000010000100000000";
-- Data_Rom(59) <= "11001001110000000000000";
-- Data_Rom(60) <= "10100000000000000000000";
-- Data_Rom(61) <= "10100000000000000000000";
-- Data_Rom(62) <= "11101000001000110000000";
-- Data_Rom(63) <= "11000000010000000000000";
-- Data_Rom(64) <= "10100000000000000000000";
-- Data_Rom(65) <= "10100000000000000000000";
-- Data_Rom(66) <= "01111010000000000000000";
-- Data_Rom(67) <= "11000110101000000000000";
-- Data_Rom(68) <= "10100000000000000000000";
-- Data_Rom(69) <= "10100000000000000000000";
-- Data_Rom(70) <= "01001000010000100000000";
-- Data_Rom(71) <= "11001000110000000000000";
-- Data_Rom(72) <= "10100000000000000000000";
-- Data_Rom(73) <= "10100000000000000000000";
-- Data_Rom(74) <= "01111010000000000000000";
-- Data_Rom(75) <= "11000111010000000000000";
-- Data_Rom(76) <= "10100000000000000000000";
-- Data_Rom(77) <= "10100000000000000000000";
-- Data_Rom(78) <= "00100010001000010000000";
-- Data_Rom(79) <= "01111010000000000000000";
-- Data_Rom(80) <= "11000111110000000000000";
-- Data_Rom(81) <= "10100000000000000000000";
-- Data_Rom(82) <= "10100000000000000000000";
-- Data_Rom(83) <= "10001000010000100000000";
-- Data_Rom(84) <= "11001010011000000000000";
-- Data_Rom(85) <= "10100000000000000000000";
-- Data_Rom(86) <= "10100000000000000000000";
-- Data_Rom(87) <= "00100010001000010000000";
-- Data_Rom(88) <= "01111010000000000000000";
-- Data_Rom(89) <= "11000000010000000000000";
-- Data_Rom(90) <= "10100000000000000000000";
-- Data_Rom(91) <= "10100000000000000000000";










-- rw='1' alors lecture
	acces_rom:process(clk)
		begin
		
		if rising_edge(clk) then
			if en='1'then
				Data_out <= Data_Rom(to_integer(unsigned(Address)));
			end if;

		end if;	
		
	end process acces_rom;

end rom_a;
