library ieee;

use IEEE.STD_LOGIC_1164.ALL;
Use ieee.numeric_std.all ;
use std.standard.all ;


entity rom is
	port(
			en			:	in std_logic;
			clk		:	in std_logic;
			Address	:	in std_logic_vector(31 downto 0);
			Data_out:	out std_logic_vector(31 downto 0)
			);
end rom;

architecture rom_a of rom is

type rom is array(0 to 4096) of std_logic_vector(7 downto 0);

signal Data_Rom : rom ;
signal Address_int : integer;
	


--------------- BEGIN -----------------------------------------------------------------
begin

Address_int <= to_integer(unsigned(Address(11 downto 0)));

-- Code here

Data_Rom(0) <= "00010011";
Data_Rom(1) <= "00000000";
Data_Rom(2) <= "00000000";
Data_Rom(3) <= "00000000";
Data_Rom(4) <= "00010011";
Data_Rom(5) <= "00000000";
Data_Rom(6) <= "00000000";
Data_Rom(7) <= "00000000";
Data_Rom(8) <= "00010011";
Data_Rom(9) <= "00000001";
Data_Rom(10) <= "00000000";
Data_Rom(11) <= "01111101";
Data_Rom(12) <= "11101111";
Data_Rom(13) <= "00000000";
Data_Rom(14) <= "10000000";
Data_Rom(15) <= "00000001";
Data_Rom(16) <= "00010011";
Data_Rom(17) <= "00000000";
Data_Rom(18) <= "00000000";
Data_Rom(19) <= "00000000";
Data_Rom(20) <= "00010011";
Data_Rom(21) <= "00000000";
Data_Rom(22) <= "00000000";
Data_Rom(23) <= "00000000";
Data_Rom(24) <= "00010011";
Data_Rom(25) <= "00000000";
Data_Rom(26) <= "00000000";
Data_Rom(27) <= "00000000";
Data_Rom(28) <= "00010011";
Data_Rom(29) <= "00000000";
Data_Rom(30) <= "00000000";
Data_Rom(31) <= "00000000";
Data_Rom(32) <= "11101111";
Data_Rom(33) <= "11110000";
Data_Rom(34) <= "10011111";
Data_Rom(35) <= "11111111";
Data_Rom(36) <= "00010011";
Data_Rom(37) <= "00000000";
Data_Rom(38) <= "00000000";
Data_Rom(39) <= "00000000";
Data_Rom(40) <= "00010011";
Data_Rom(41) <= "00000001";
Data_Rom(42) <= "11000001";
Data_Rom(43) <= "11111111";
Data_Rom(44) <= "00100011";
Data_Rom(45) <= "00100000";
Data_Rom(46) <= "00010001";
Data_Rom(47) <= "00000000";
Data_Rom(48) <= "00010011";
Data_Rom(49) <= "00000001";
Data_Rom(50) <= "11000001";
Data_Rom(51) <= "11111111";
Data_Rom(52) <= "10010011";
Data_Rom(53) <= "00000110";
Data_Rom(54) <= "00000000";
Data_Rom(55) <= "00000000";
Data_Rom(56) <= "00010011";
Data_Rom(57) <= "00000110";
Data_Rom(58) <= "00000000";
Data_Rom(59) <= "00000000";
Data_Rom(60) <= "00110011";
Data_Rom(61) <= "00000110";
Data_Rom(62) <= "11010110";
Data_Rom(63) <= "00000000";
Data_Rom(64) <= "00110011";
Data_Rom(65) <= "00000110";
Data_Rom(66) <= "11010110";
Data_Rom(67) <= "00000000";
Data_Rom(68) <= "00110011";
Data_Rom(69) <= "00000110";
Data_Rom(70) <= "11010110";
Data_Rom(71) <= "00000000";
Data_Rom(72) <= "00110011";
Data_Rom(73) <= "00000110";
Data_Rom(74) <= "11010110";
Data_Rom(75) <= "00000000";
Data_Rom(76) <= "10010111";
Data_Rom(77) <= "00000010";
Data_Rom(78) <= "00000000";
Data_Rom(79) <= "00000000";
Data_Rom(80) <= "10010011";
Data_Rom(81) <= "10000010";
Data_Rom(82) <= "11000010";
Data_Rom(83) <= "00000000";
Data_Rom(84) <= "00110011";
Data_Rom(85) <= "00000110";
Data_Rom(86) <= "01010110";
Data_Rom(87) <= "00000000";
Data_Rom(88) <= "00000011";
Data_Rom(89) <= "00101111";
Data_Rom(90) <= "01000110";
Data_Rom(91) <= "00011011";
Data_Rom(92) <= "10010011";
Data_Rom(93) <= "00000011";
Data_Rom(94) <= "00010000";
Data_Rom(95) <= "00000000";
Data_Rom(96) <= "00010011";
Data_Rom(97) <= "00000011";
Data_Rom(98) <= "00000000";
Data_Rom(99) <= "00000000";
Data_Rom(100) <= "00110011";
Data_Rom(101) <= "00000011";
Data_Rom(102) <= "11010011";
Data_Rom(103) <= "00000000";
Data_Rom(104) <= "00110011";
Data_Rom(105) <= "00000011";
Data_Rom(106) <= "11010011";
Data_Rom(107) <= "00000000";
Data_Rom(108) <= "00110011";
Data_Rom(109) <= "00000011";
Data_Rom(110) <= "11010011";
Data_Rom(111) <= "00000000";
Data_Rom(112) <= "00110011";
Data_Rom(113) <= "00000011";
Data_Rom(114) <= "11010011";
Data_Rom(115) <= "00000000";
Data_Rom(116) <= "10010111";
Data_Rom(117) <= "00000010";
Data_Rom(118) <= "00000000";
Data_Rom(119) <= "00000000";
Data_Rom(120) <= "10010011";
Data_Rom(121) <= "10000010";
Data_Rom(122) <= "11000010";
Data_Rom(123) <= "00000000";
Data_Rom(124) <= "00110011";
Data_Rom(125) <= "00000011";
Data_Rom(126) <= "01010011";
Data_Rom(127) <= "00000000";
Data_Rom(128) <= "00100011";
Data_Rom(129) <= "00100110";
Data_Rom(130) <= "01110011";
Data_Rom(131) <= "00011000";
Data_Rom(132) <= "10010011";
Data_Rom(133) <= "00001111";
Data_Rom(134) <= "00010000";
Data_Rom(135) <= "00000000";
Data_Rom(136) <= "00010011";
Data_Rom(137) <= "00001110";
Data_Rom(138) <= "00000000";
Data_Rom(139) <= "00000000";
Data_Rom(140) <= "00110011";
Data_Rom(141) <= "00001110";
Data_Rom(142) <= "11111110";
Data_Rom(143) <= "00000001";
Data_Rom(144) <= "00110011";
Data_Rom(145) <= "00001110";
Data_Rom(146) <= "11111110";
Data_Rom(147) <= "00000001";
Data_Rom(148) <= "00110011";
Data_Rom(149) <= "00001110";
Data_Rom(150) <= "11111110";
Data_Rom(151) <= "00000001";
Data_Rom(152) <= "00110011";
Data_Rom(153) <= "00001110";
Data_Rom(154) <= "11111110";
Data_Rom(155) <= "00000001";
Data_Rom(156) <= "10010111";
Data_Rom(157) <= "00000010";
Data_Rom(158) <= "00000000";
Data_Rom(159) <= "00000000";
Data_Rom(160) <= "10010011";
Data_Rom(161) <= "10000010";
Data_Rom(162) <= "11000010";
Data_Rom(163) <= "00000000";
Data_Rom(164) <= "00110011";
Data_Rom(165) <= "00001110";
Data_Rom(166) <= "01011110";
Data_Rom(167) <= "00000000";
Data_Rom(168) <= "10000011";
Data_Rom(169) <= "00100010";
Data_Rom(170) <= "01001110";
Data_Rom(171) <= "00010110";
Data_Rom(172) <= "10010011";
Data_Rom(173) <= "00000011";
Data_Rom(174) <= "00010000";
Data_Rom(175) <= "00000000";
Data_Rom(176) <= "00010011";
Data_Rom(177) <= "00000011";
Data_Rom(178) <= "00000000";
Data_Rom(179) <= "00000000";
Data_Rom(180) <= "00110011";
Data_Rom(181) <= "00000011";
Data_Rom(182) <= "11110011";
Data_Rom(183) <= "00000001";
Data_Rom(184) <= "00110011";
Data_Rom(185) <= "00000011";
Data_Rom(186) <= "11110011";
Data_Rom(187) <= "00000001";
Data_Rom(188) <= "00110011";
Data_Rom(189) <= "00000011";
Data_Rom(190) <= "11110011";
Data_Rom(191) <= "00000001";
Data_Rom(192) <= "00110011";
Data_Rom(193) <= "00000011";
Data_Rom(194) <= "11110011";
Data_Rom(195) <= "00000001";
Data_Rom(196) <= "10010111";
Data_Rom(197) <= "00000010";
Data_Rom(198) <= "00000000";
Data_Rom(199) <= "00000000";
Data_Rom(200) <= "10010011";
Data_Rom(201) <= "10000010";
Data_Rom(202) <= "11000010";
Data_Rom(203) <= "00000000";
Data_Rom(204) <= "00110011";
Data_Rom(205) <= "00000011";
Data_Rom(206) <= "01010011";
Data_Rom(207) <= "00000000";
Data_Rom(208) <= "00100011";
Data_Rom(209) <= "00101110";
Data_Rom(210) <= "01110011";
Data_Rom(211) <= "00010010";
Data_Rom(212) <= "10000011";
Data_Rom(213) <= "00100010";
Data_Rom(214) <= "00000001";
Data_Rom(215) <= "00000000";
Data_Rom(216) <= "10010011";
Data_Rom(217) <= "00000010";
Data_Rom(218) <= "00100000";
Data_Rom(219) <= "00000000";
Data_Rom(220) <= "00100011";
Data_Rom(221) <= "00100000";
Data_Rom(222) <= "01010001";
Data_Rom(223) <= "00000000";
Data_Rom(224) <= "00010011";
Data_Rom(225) <= "00000000";
Data_Rom(226) <= "00000000";
Data_Rom(227) <= "00000000";
Data_Rom(228) <= "10000011";
Data_Rom(229) <= "00100011";
Data_Rom(230) <= "00000001";
Data_Rom(231) <= "00000000";
Data_Rom(232) <= "00010011";
Data_Rom(233) <= "00000011";
Data_Rom(234) <= "10000000";
Data_Rom(235) <= "00000000";
Data_Rom(236) <= "10110011";
Data_Rom(237) <= "10000010";
Data_Rom(238) <= "01100011";
Data_Rom(239) <= "01000000";
Data_Rom(240) <= "01100011";
Data_Rom(241) <= "11000110";
Data_Rom(242) <= "00000010";
Data_Rom(243) <= "00000000";
Data_Rom(244) <= "10010011";
Data_Rom(245) <= "00000010";
Data_Rom(246) <= "00010000";
Data_Rom(247) <= "00000000";
Data_Rom(248) <= "11101111";
Data_Rom(249) <= "00000000";
Data_Rom(250) <= "10000000";
Data_Rom(251) <= "00000000";
Data_Rom(252) <= "10010011";
Data_Rom(253) <= "00000010";
Data_Rom(254) <= "00000000";
Data_Rom(255) <= "00000000";
Data_Rom(256) <= "01100011";
Data_Rom(257) <= "10010110";
Data_Rom(258) <= "00000010";
Data_Rom(259) <= "00001100";
Data_Rom(260) <= "10000011";
Data_Rom(261) <= "00101110";
Data_Rom(262) <= "00000001";
Data_Rom(263) <= "00000000";
Data_Rom(264) <= "00010011";
Data_Rom(265) <= "00000011";
Data_Rom(266) <= "00000000";
Data_Rom(267) <= "00000000";
Data_Rom(268) <= "00110011";
Data_Rom(269) <= "00000011";
Data_Rom(270) <= "11010011";
Data_Rom(271) <= "00000001";
Data_Rom(272) <= "00110011";
Data_Rom(273) <= "00000011";
Data_Rom(274) <= "11010011";
Data_Rom(275) <= "00000001";
Data_Rom(276) <= "00110011";
Data_Rom(277) <= "00000011";
Data_Rom(278) <= "11010011";
Data_Rom(279) <= "00000001";
Data_Rom(280) <= "00110011";
Data_Rom(281) <= "00000011";
Data_Rom(282) <= "11010011";
Data_Rom(283) <= "00000001";
Data_Rom(284) <= "10010111";
Data_Rom(285) <= "00000010";
Data_Rom(286) <= "00000000";
Data_Rom(287) <= "00000000";
Data_Rom(288) <= "10010011";
Data_Rom(289) <= "10000010";
Data_Rom(290) <= "11000010";
Data_Rom(291) <= "00000000";
Data_Rom(292) <= "00110011";
Data_Rom(293) <= "00000011";
Data_Rom(294) <= "01010011";
Data_Rom(295) <= "00000000";
Data_Rom(296) <= "10000011";
Data_Rom(297) <= "00100010";
Data_Rom(298) <= "01000011";
Data_Rom(299) <= "00001110";
Data_Rom(300) <= "00000011";
Data_Rom(301) <= "00100011";
Data_Rom(302) <= "00000001";
Data_Rom(303) <= "00000000";
Data_Rom(304) <= "10010011";
Data_Rom(305) <= "00000010";
Data_Rom(306) <= "00100000";
Data_Rom(307) <= "00000000";
Data_Rom(308) <= "10110011";
Data_Rom(309) <= "00000011";
Data_Rom(310) <= "01010011";
Data_Rom(311) <= "01000000";
Data_Rom(312) <= "00010011";
Data_Rom(313) <= "00000011";
Data_Rom(314) <= "00000000";
Data_Rom(315) <= "00000000";
Data_Rom(316) <= "00110011";
Data_Rom(317) <= "00000011";
Data_Rom(318) <= "01110011";
Data_Rom(319) <= "00000000";
Data_Rom(320) <= "00110011";
Data_Rom(321) <= "00000011";
Data_Rom(322) <= "01110011";
Data_Rom(323) <= "00000000";
Data_Rom(324) <= "00110011";
Data_Rom(325) <= "00000011";
Data_Rom(326) <= "01110011";
Data_Rom(327) <= "00000000";
Data_Rom(328) <= "00110011";
Data_Rom(329) <= "00000011";
Data_Rom(330) <= "01110011";
Data_Rom(331) <= "00000000";
Data_Rom(332) <= "10010111";
Data_Rom(333) <= "00000010";
Data_Rom(334) <= "00000000";
Data_Rom(335) <= "00000000";
Data_Rom(336) <= "10010011";
Data_Rom(337) <= "10000010";
Data_Rom(338) <= "11000010";
Data_Rom(339) <= "00000000";
Data_Rom(340) <= "00110011";
Data_Rom(341) <= "00000011";
Data_Rom(342) <= "01010011";
Data_Rom(343) <= "00000000";
Data_Rom(344) <= "00000011";
Data_Rom(345) <= "00101110";
Data_Rom(346) <= "01000011";
Data_Rom(347) <= "00001011";
Data_Rom(348) <= "00000011";
Data_Rom(349) <= "00100011";
Data_Rom(350) <= "00000001";
Data_Rom(351) <= "00000000";
Data_Rom(352) <= "10010011";
Data_Rom(353) <= "00000010";
Data_Rom(354) <= "00010000";
Data_Rom(355) <= "00000000";
Data_Rom(356) <= "10110011";
Data_Rom(357) <= "00000011";
Data_Rom(358) <= "01010011";
Data_Rom(359) <= "01000000";
Data_Rom(360) <= "00010011";
Data_Rom(361) <= "00000011";
Data_Rom(362) <= "00000000";
Data_Rom(363) <= "00000000";
Data_Rom(364) <= "00110011";
Data_Rom(365) <= "00000011";
Data_Rom(366) <= "01110011";
Data_Rom(367) <= "00000000";
Data_Rom(368) <= "00110011";
Data_Rom(369) <= "00000011";
Data_Rom(370) <= "01110011";
Data_Rom(371) <= "00000000";
Data_Rom(372) <= "00110011";
Data_Rom(373) <= "00000011";
Data_Rom(374) <= "01110011";
Data_Rom(375) <= "00000000";
Data_Rom(376) <= "00110011";
Data_Rom(377) <= "00000011";
Data_Rom(378) <= "01110011";
Data_Rom(379) <= "00000000";
Data_Rom(380) <= "10010111";
Data_Rom(381) <= "00000010";
Data_Rom(382) <= "00000000";
Data_Rom(383) <= "00000000";
Data_Rom(384) <= "10010011";
Data_Rom(385) <= "10000010";
Data_Rom(386) <= "11000010";
Data_Rom(387) <= "00000000";
Data_Rom(388) <= "00110011";
Data_Rom(389) <= "00000011";
Data_Rom(390) <= "01010011";
Data_Rom(391) <= "00000000";
Data_Rom(392) <= "10000011";
Data_Rom(393) <= "00100010";
Data_Rom(394) <= "01000011";
Data_Rom(395) <= "00001000";
Data_Rom(396) <= "10110011";
Data_Rom(397) <= "00000011";
Data_Rom(398) <= "01011110";
Data_Rom(399) <= "00000000";
Data_Rom(400) <= "00010011";
Data_Rom(401) <= "00000011";
Data_Rom(402) <= "00000000";
Data_Rom(403) <= "00000000";
Data_Rom(404) <= "00110011";
Data_Rom(405) <= "00000011";
Data_Rom(406) <= "11010011";
Data_Rom(407) <= "00000001";
Data_Rom(408) <= "00110011";
Data_Rom(409) <= "00000011";
Data_Rom(410) <= "11010011";
Data_Rom(411) <= "00000001";
Data_Rom(412) <= "00110011";
Data_Rom(413) <= "00000011";
Data_Rom(414) <= "11010011";
Data_Rom(415) <= "00000001";
Data_Rom(416) <= "00110011";
Data_Rom(417) <= "00000011";
Data_Rom(418) <= "11010011";
Data_Rom(419) <= "00000001";
Data_Rom(420) <= "10010111";
Data_Rom(421) <= "00000010";
Data_Rom(422) <= "00000000";
Data_Rom(423) <= "00000000";
Data_Rom(424) <= "10010011";
Data_Rom(425) <= "10000010";
Data_Rom(426) <= "11000010";
Data_Rom(427) <= "00000000";
Data_Rom(428) <= "00110011";
Data_Rom(429) <= "00000011";
Data_Rom(430) <= "01010011";
Data_Rom(431) <= "00000000";
Data_Rom(432) <= "00100011";
Data_Rom(433) <= "00101110";
Data_Rom(434) <= "01110011";
Data_Rom(435) <= "00000100";
Data_Rom(436) <= "10000011";
Data_Rom(437) <= "00100010";
Data_Rom(438) <= "00000001";
Data_Rom(439) <= "00000000";
Data_Rom(440) <= "10000011";
Data_Rom(441) <= "00100011";
Data_Rom(442) <= "00000001";
Data_Rom(443) <= "00000000";
Data_Rom(444) <= "00010011";
Data_Rom(445) <= "00000011";
Data_Rom(446) <= "00010000";
Data_Rom(447) <= "00000000";
Data_Rom(448) <= "10110011";
Data_Rom(449) <= "10000010";
Data_Rom(450) <= "01100011";
Data_Rom(451) <= "00000000";
Data_Rom(452) <= "00100011";
Data_Rom(453) <= "00100000";
Data_Rom(454) <= "01010001";
Data_Rom(455) <= "00000000";
Data_Rom(456) <= "11101111";
Data_Rom(457) <= "11110000";
Data_Rom(458) <= "10011111";
Data_Rom(459) <= "11110001";
Data_Rom(460) <= "10010011";
Data_Rom(461) <= "00000010";
Data_Rom(462) <= "01110000";
Data_Rom(463) <= "00000000";
Data_Rom(464) <= "00010011";
Data_Rom(465) <= "00000011";
Data_Rom(466) <= "00000000";
Data_Rom(467) <= "00000000";
Data_Rom(468) <= "00110011";
Data_Rom(469) <= "00000011";
Data_Rom(470) <= "01010011";
Data_Rom(471) <= "00000000";
Data_Rom(472) <= "00110011";
Data_Rom(473) <= "00000011";
Data_Rom(474) <= "01010011";
Data_Rom(475) <= "00000000";
Data_Rom(476) <= "00110011";
Data_Rom(477) <= "00000011";
Data_Rom(478) <= "01010011";
Data_Rom(479) <= "00000000";
Data_Rom(480) <= "00110011";
Data_Rom(481) <= "00000011";
Data_Rom(482) <= "01010011";
Data_Rom(483) <= "00000000";
Data_Rom(484) <= "10010111";
Data_Rom(485) <= "00000010";
Data_Rom(486) <= "00000000";
Data_Rom(487) <= "00000000";
Data_Rom(488) <= "10010011";
Data_Rom(489) <= "10000010";
Data_Rom(490) <= "11000010";
Data_Rom(491) <= "00000000";
Data_Rom(492) <= "00110011";
Data_Rom(493) <= "00000011";
Data_Rom(494) <= "01010011";
Data_Rom(495) <= "00000000";
Data_Rom(496) <= "10000011";
Data_Rom(497) <= "00100010";
Data_Rom(498) <= "11000011";
Data_Rom(499) <= "00000001";
Data_Rom(500) <= "00010011";
Data_Rom(501) <= "10000101";
Data_Rom(502) <= "00000010";
Data_Rom(503) <= "00000000";
Data_Rom(504) <= "11101111";
Data_Rom(505) <= "00000000";
Data_Rom(506) <= "01000000";
Data_Rom(507) <= "00000000";
Data_Rom(508) <= "00010011";
Data_Rom(509) <= "00000000";
Data_Rom(510) <= "00000000";
Data_Rom(511) <= "00000000";
Data_Rom(512) <= "10000011";
Data_Rom(513) <= "00100000";
Data_Rom(514) <= "01000001";
Data_Rom(515) <= "00000000";
Data_Rom(516) <= "00010011";
Data_Rom(517) <= "00000001";
Data_Rom(518) <= "11000001";
Data_Rom(519) <= "00000000";
Data_Rom(520) <= "11100111";
Data_Rom(521) <= "10000000";
Data_Rom(522) <= "00000000";
Data_Rom(523) <= "00000000";


	acces_rom:process(clk)
		begin
		
		if rising_edge(clk) then
			if en='1'then
				Data_out <= Data_Rom(Address_int+3) & Data_Rom(Address_int+2) &
							Data_Rom(Address_int+1) & Data_Rom(Address_int);
			end if;

		end if;	
		
	end process acces_rom;

end rom_a;
